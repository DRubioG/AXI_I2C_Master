
--! Registros
--! ==
--! | Nombre  | Offset | R/W | Descripci�n |
--! |---------|--------|-----|-------------|
--! | CNTRL   |   0x0  |  W  | Registro de control del bloque IP |
--! | WRITE   |   0x4  |  W  | Registro para escribir por I2C |
--! | READ    |   0x8  |  R  | Registro para leer por I2C |
--!
--! CNTRL
--! --
--! - **EN**: Bit de habilitaci�n del bloque IP.
--! - **ST**: Bit de start de la interfaz I2C.
--! - **SP**: Bit de parada de la interfaz I2C.
--! - **RD**: Bit de lectura de la interfaz I2C.
--! - **FF**: Bit de lectura del FIFO
--! {
--!       "config": { 
--!         "hspace": 1000
--!       },
--!     reg:[
--!     { "name": "EN",   		"bits": 1, "attr": "w", "type": 4},
--!     { "name": "ST",   		"bits": 1, "attr": "w", "type": 5 },
--!     { "name": "SP",   		"bits": 1, "attr": "w", "type": 6 },
--!     { "name": "RD",   		"bits": 1, "attr": "w", "type": 7 },
--!     { "name": "FF",   		"bits": 1, "attr": "w", "type": 2 },
--!     { "name": "Size",   	"bits": 8, "attr": "w", "type": 3 },
--!     { "name": "Reserved",   "bits": 19, "attr": "", "type":"not used" }
--! ]}
--! WRITE
--! --
--! - **Address**: Direcci�n de escritura del I2C.
--! - **Data**: Dato a escribir por I2C.
--! {
--!       "config": { 
--!         "hspace": 1000
--!       },
--!     reg:[
--!     { "name": "Address",   	"bits": 7, "attr": "w", "type":2 },
--!     { "name": "Data",   	"bits": 8, "attr": "w", "type":3 },
--!     { "name": "Reserved",   "bits": 17, "attr": "", "type":"not used" }
--! ]}
--! READ
--! --
--! - **Data**: Dato le�do por I2C.
--! {
--!       "config": { 
--!         "hspace": 1000
--!       },
--!     reg:[
--!     { "name": "Data",   	"bits": 8, "attr": "r" , "type": 4},
--!     { "name": "Reserved",   "bits": 24, "attr": "", "type":"not used" }
--! ]}

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity AXI_I2C_Master is
	generic (
		-- Users to add parameters here

		-- User parameters ends
		-- Do not modify the parameters beyond this line


		-- Parameters of Axi Slave Bus Interface S_AXI
		C_S_AXI_DATA_WIDTH	: integer	:= 32;
		C_S_AXI_ADDR_WIDTH	: integer	:= 4
	);
	port (
		-- Users to add ports here
		SDA : inout std_logic;
		SCL : out std_logic;
		-- User ports ends
		-- Do not modify the ports beyond this line


		-- Ports of Axi Slave Bus Interface S_AXI
		--! @virtualbus AXI @dir in
		s_axi_aclk	: in std_logic;
		s_axi_aresetn	: in std_logic;
		s_axi_awaddr	: in std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
		s_axi_awprot	: in std_logic_vector(2 downto 0);
		s_axi_awvalid	: in std_logic;
		s_axi_awready	: out std_logic;
		s_axi_wdata	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
		s_axi_wstrb	: in std_logic_vector((C_S_AXI_DATA_WIDTH/8)-1 downto 0);
		s_axi_wvalid	: in std_logic;
		s_axi_wready	: out std_logic;
		s_axi_bresp	: out std_logic_vector(1 downto 0);
		s_axi_bvalid	: out std_logic;
		s_axi_bready	: in std_logic;
		s_axi_araddr	: in std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
		s_axi_arprot	: in std_logic_vector(2 downto 0);
		s_axi_arvalid	: in std_logic;
		s_axi_arready	: out std_logic;
		s_axi_rdata	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
		s_axi_rresp	: out std_logic_vector(1 downto 0);
		s_axi_rvalid	: out std_logic;
		s_axi_rready	: in std_logic
		--! @end
	);
end AXI_I2C_Master;

architecture arch_imp of AXI_I2C_Master is

begin

-- Instantiation of Axi Bus Interface S_AXI
AXI_I2C_Master_slave_lite_v1_0_S_AXI_inst : entity work.AXI_I2C_Master_slave_lite_v1_0_S_AXI
	generic map (
		C_S_AXI_DATA_WIDTH	=> C_S_AXI_DATA_WIDTH,
		C_S_AXI_ADDR_WIDTH	=> C_S_AXI_ADDR_WIDTH
	)
	port map (
		SDA => SDA,
		SCL => SCL,
		S_AXI_ACLK	=> s_axi_aclk,
		S_AXI_ARESETN	=> s_axi_aresetn,
		S_AXI_AWADDR	=> s_axi_awaddr,
		S_AXI_AWPROT	=> s_axi_awprot,
		S_AXI_AWVALID	=> s_axi_awvalid,
		S_AXI_AWREADY	=> s_axi_awready,
		S_AXI_WDATA	=> s_axi_wdata,
		S_AXI_WSTRB	=> s_axi_wstrb,
		S_AXI_WVALID	=> s_axi_wvalid,
		S_AXI_WREADY	=> s_axi_wready,
		S_AXI_BRESP	=> s_axi_bresp,
		S_AXI_BVALID	=> s_axi_bvalid,
		S_AXI_BREADY	=> s_axi_bready,
		S_AXI_ARADDR	=> s_axi_araddr,
		S_AXI_ARPROT	=> s_axi_arprot,
		S_AXI_ARVALID	=> s_axi_arvalid,
		S_AXI_ARREADY	=> s_axi_arready,
		S_AXI_RDATA	=> s_axi_rdata,
		S_AXI_RRESP	=> s_axi_rresp,
		S_AXI_RVALID	=> s_axi_rvalid,
		S_AXI_RREADY	=> s_axi_rready
	);

	-- Add user logic here

	-- User logic ends

end arch_imp;
